{"api/toc.html":"314rtfz3.kvq","articles/toc.html":"lposw313.pam","ProcessDoku/SalesProcess copy 2.html":"sooherin.wju","ProcessDoku/toc.html":"yr3gtopp.3mx","toc.html":"fi0qkohp.zk0","ProcessDoku/intro.html":"lvhoyazj.om2","articles/SalesProcess.html":"i4d3o43s.0xw","ProcessDoku/SalesProcess copy 5.html":"rmj2uydg.rso","ProcessDoku/SalesProcess copy 4.html":"j55kj5r5.so5","ProcessDoku/SalesProcess copy 3.html":"uc2ibhhj.g42","api/index.html":"ky43qtut.lxa","ProcessDoku/SalesProcess copy 6.html":"e4mtvijm.pm5","api/index1.html":"c1yfevou.spo","index.html":"atmmo1pf.3o4","ProcessDoku/SalesProcess.html":"dxmhwt34.zva","ProcessDoku/SalesProcess copy 7.html":"vyplwhtv.2gm","articles/intro.html":"h54jkbrn.clb","ProcessDoku/SalesProcess copy.html":"v22is5fm.0cw"}