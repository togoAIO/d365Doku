<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Neuigkeiten oder &#196;nderungen in Dynamics 365 Talent (30. April, 2019) | WIKA Documentation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Neuigkeiten oder &#196;nderungen in Dynamics 365 Talent (30. April, 2019) | WIKA Documentation ">
    <meta name="generator" content="docfx 2.56.6.0">
    
    <link rel="shortcut icon" href="../../microsoft-dynamics-crm-365-icon.ico">
    <link rel="stylesheet" href="../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../styles/docfx.css">
    <link rel="stylesheet" href="../../styles/main.css">
    <link href="https://fonts.googleapis.com/css?family=Roboto" rel="stylesheet"> 
    <meta property="docfx:navrel" content="../../toc.html">
    <meta property="docfx:tocrel" content="TOC.html">
    
    
    
  </head>  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../index.html">
                <img id="logo" class="svg" src="../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="">
<h1 id="whats-new-or-changed-in-dynamics-365-talent-april-30-2019" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="28">Neuigkeiten oder Änderungen in Dynamics 365 Talent (30. April, 2019)</h1>

[!include[rename-banner](~/includes/cc-data-platform-banner.md)]
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="32">In diesem Thema werden die Funktionen beschrieben, die in Microsoft Dynamics 365 Talent entweder neu oder geändert sind.</p>
<h2 id="changes-in-attract" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="34">Änderungen in Attract</h2>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="36">Diese Version enthält kleinere Fehlerkorrekturen für Dynamics 365 Talent: Attract.</p>
<h2 id="changes-in-onboard" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="38">Änderungen in Onboard</h2>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="40">Diese Version enthält kleinere Fehlerkorrekturen für Dynamics 365 Talent: Onboard.</p>
<h2 id="changes-in-core-hr" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="42">Core HR-Änderungen</h2>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="44">Die in diesem Abschnitt beschriebenen Änderungen gelten für Buildnummer 8.1.2270. Die Zahlen in Klammern in einigen Überschriften beziehen sich auf Supportnummern in Microsoft Dynamics Lifecycle Services (LCS).</p>
<h3 id="provide-feedback" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="46">Feedback geben</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="48">Die Option, zum Bereitstellen von Feedback befindet sich im Menü <strong sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="48">Hilfe</strong> (<strong sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="48">?</strong>) in Talent. Dieses Menü bietet Zugriff auf den folgenden Ressourcen:</p>
<ul sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="50">
<li sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="50">Feedback</li>
<li sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="51">Hilfe</li>
<li sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="52">Erste Schritte</li>
<li sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="53">Unterstützung</li>
<li sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="54">Ideen</li>
<li sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="55">Info</li>
</ul>
<h3 id="improvements-to-the-user-interface-for-duplicate-employee-detection" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="57">Verbesserungen an der Benutzeroberfläche, um doppelten Mitarbeiter zu erkennen</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="59">Aufgrund dieser Änderung werden Duplikate nun beim Festlegen von Namensfeldern erkannt und eine Statusanzeige zeigt die Anzahl der Duplikate an, die erfasst wurden. Ein bereitgestellter Link öffnet eine Seite, auf der Sie bewerten können, ob Sie eines der Duplikate verwenden sollen. Die Duplikatsseite wird nicht automatisch geöffnet, damit die Dateneingabe nicht unterbrochen wird. Sie müssen den Link auswählen, um die Seite zu öffnen.</p>
<h3 id="common-data-service-entity-support-for-custom-fields" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="61">Common Data Service-Entitätssupport für benutzerdefinierte Felder</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="63">In der Version dieser Woche unterstützen die folgenden Entitäten nun benutzerdefinierte Felder: Anstellung, Vorteilstyp und Lohnzyklus.</p>
<h3 id="an-error-occurs-when-an-off-boarding-checklist-is-assigned-299877" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="65">Ein Fehler tritt auf, wenn eine Offboarding-Checkliste zugeordnet wird (299877 )</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="67">Mit dieser Änderung wird eine Fehlermeldung korrigiert, die angezeigt wird, wenn Sie einem Mitarbeiter außerhalb des Kündigungsprozesses eine Offboarding-Checkliste zuweisen.</p>
<h3 id="the-exited-workers-link-opens-the-wrong-worker-309939" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="69">Der Link für beendete Arbeitskräfte öffnet die falsche Arbeitskraft (309939)</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="71">Mit dieser Änderung wird ein Problem behoben, das auftritt, wenn Sie einen Mitarbeiter aus einer anderen juristischen Person neu anwerben und versuchen, aus der Liste der beendeten Arbeitskräfte zu dem Mitarbeiter zu wechseln.</p>
<h3 id="the-employee-self-service-compensation-card-doesnt-show-summary-values-when-advanced-security-is-turned-on-315231" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="73">Die Mitarbeiter-Self-Service-Kompensationskarte zeigt keine Zusammenfassungswerte an, wenn die erweiterte Sicherheit eingeschaltet wird (315231 )</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="75">Mit dieser Änderung wird ein Problem behoben, das auftritt, wenn Sie erweiterte Kompensationssicherheit verwenden. Wenn die erweiterte Sicherheit aktiviert ist, zeigt der Mitarbeiter-Self-Service nun die zusammengefassten Kompensationsbeträge für Mitarbeiter und Manager an. Vor dieser Änderung wurden zusammenfassende Werte als 0 (null) angezeigt.</p>
<h3 id="if-a-position-without-a-title-is-created-in-common-data-service-no-position-is-created-in-talent-314562" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="77">Wenn eine Position ohne einen Titel in Common Data Service erstellt wird, wird keine Position im Talent erstellt(314562)</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="79">Mit den Änderungen dieser Woche wird ein Problem behoben, das auftritt, wenn Sie Positionen in Common Data Service erstellen, jedoch keinen Titel hinzufügen.</p>
<h3 id="error-message-in-performance-journal-entries-in-employee-self-service-314134" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="81">Fehlermeldung in den Leistungsjournaleinträgen im Mitarbeiter-Self-Service (314134 )</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="83">Mit dieser Änderung wird ein Problem behoben, das auftritt, wenn Sie den Leistungsjournaleinträgen Leistungsziele im Mitarbeiter-Self-Service zuordnen.</p>
<h2 id="in-preview" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="85">Vorschau</h2>
<h3 id="allow-reason-codes-to-be-specified-on-leave-types" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="87">Ermöglichen Sie, dass Ursachencodes für Sonderurlaubstypen angegeben werden können</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="89">Organisationen brauchen möglicherweise zusätzliche Informationen zu Freizeitanforderungen. Sie können nun Ursachencodes für Sonderurlaubstypen definieren und Mitarbeiter aktivieren, damit sie einen Ursachencode für ihre Freizeitanforderungen auszuwählen können.</p>
<h3 id="require-reason-codes-for-specific-leave-types-on-time-off-requests" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="91">Erfordert Ursachencodes für bestimmte Urlaubstypen bei Freizeitanforderungen</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="93">Organisationen brauchen ggf. bestimmte Ursachencodes für Sonderurlaubstypen, wenn Mitarbeiter Freizeit beantragen. Diese Anforderung ist möglicherweise aufgrund der Unternehmensrichtlinie oder der gesetzlichen Vorgaben vorhanden. Sie können nun angeben, welche Urlaubstypen einen Ursachencodes erfordern und Sie können von Mitarbeitern verlangen, dass sie einen Ursachencode für den Sonderurlaubstyp für ihre Freizeitanforderungen angeben.</p>
<h3 id="provide-a-leave-and-absence-transaction-list-for-hr" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="95">Erstellen Sie eine Urlaub- und Abwesenheitsbuchungsliste für die Personalverwaltung</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="97">Die Möglichkeit zum Nachverfolgen von Mitarbeiterfreizeit und ein Verständnis dafür, wie Freizeit berechnet wird, hilft nicht nur der Personalverwaltung, Fragen von Mitarbeitern zu beantworten sondern garantiert auch, dass die Freizeit für Mitarbeiter korrekt ist. Personalverwaltung besitzt nun eine neue Anzeige in den Transaktionen (Abgrenzungen, Zuschüsse, Regulierungen und Anforderungen), sodass die Mitarbeiter der Personalverwaltung die Gründe hinter den Salden anzeigen können.</p>
<h2 id="coming-soon" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="99">Bald verfügbar</h2>
<h3 id="email-support-for-alerts" sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="101">E-Mail-Support für Warnungen</h3>
<p sourcefile="articles_de/talent/whats-new-talent-april-30-2019.md" sourcestartlinenumber="103">Durch das Plattformupdate 26 für Finance and Operations können Benutzer Warnregeln erstellen, dass automatisch E-Mail-Benachrichtigungen an Kontakte gesendet werden, wenn dies von einem Ereignis ausgelöst wird.</p>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../styles/main.js"></script>
  </body>
</html>
