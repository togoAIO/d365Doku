<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Ausschreibungstypen und Bewertungskriterien f&#252;r Angebotsanforderungen erstellen | WIKA Documentation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Ausschreibungstypen und Bewertungskriterien f&#252;r Angebotsanforderungen erstellen | WIKA Documentation ">
    <meta name="generator" content="docfx 2.56.6.0">
    
    <link rel="shortcut icon" href="../../../../microsoft-dynamics-crm-365-icon.ico">
    <link rel="stylesheet" href="../../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../../styles/main.css">
    <link href="https://fonts.googleapis.com/css?family=Roboto" rel="stylesheet"> 
    <meta property="docfx:navrel" content="../../../../toc.html">
    <meta property="docfx:tocrel" content="../../toc.html">
    
    
    
  </head>  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../../index.html">
                <img id="logo" class="svg" src="../../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="">
<h1 id="create-solicitation-types-and-scoring-criteria-for-rfqs" sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="26">Ausschreibungstypen und Bewertungskriterien für Angebotsanforderungen erstellen</h1>

<div class="IMPORTANT" sourcefile="articles_de/supply-chain/includes/banner.md" sourcestartlinenumber="1">
<h5>Important</h5>
<p sourcefile="articles_de/supply-chain/includes/banner.md" sourcestartlinenumber="2">Dynamics 365 for Finance and Operations hat sich zu speziell entwickelten Anwendungen entwickelt, mit denen Sie bestimmte Geschäftsfunktionen verwalten können. Weitere Informationen zu diesen Änderungen finden Sie im <a href="https://go.microsoft.com/fwlink/?LinkId=866544" sourcefile="articles_de/supply-chain/includes/banner.md" sourcestartlinenumber="2">Dynamics 365-Lizenzierungshandbuch</a>.</p>
</div>

<p sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="30">Dieser Leitfaden zeigt Ihnen, wie man einen Ausschreibungstyp erstellt und diesen einer Bewertungsmethode zuordnet. Er zeigt auch, wie man den Ausschreibungstyp auf eine Angebotsanforderung anwendet, wodurch die Standardbewertungsmethode festgelegt wird. Diese Aufgaben werden normalerweise von einem Einkaufsleiter ausgeführt. Sie können diese Prozedur im Demodatenunternehmen USMF oder für Ihre eigenen Daten verwenden. Sie müssen eine Bewertungsmethode verfügbar haben, bevor Sie beginnen.</p>
<h2 id="create-a-solicitation-type" sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="33">Erstellt eines neuen Anforderungstyps</h2>
<ol sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="34">
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="34">Wechseln Sie zu Beschaffung &gt; Einstellungen &gt; Angebotsanforderung &gt; Anforderungstyp.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="35">Klicken Sie auf &quot;Neu&quot;.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="36">Geben Sie im Feld &quot;Name&quot; einen Wert ein.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="37">Geben Sie im Feld &quot;Beschreibung&quot; einen Wert ein.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="38">Wählen Sie im Feld &quot;Bewertungsmethode&quot; die Bewertungsmethode aus, die Sie für diesen Ausschreibungstyp verwenden möchten.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="39">Klicken Sie auf &quot;Speichern&quot;.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="40">Schließen Sie die Seite.</li>
</ol>
<h2 id="use-the-solicitation-type" sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="42">Den Ausschreibungstyp verwenden</h2>
<ol sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="43">
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="43">Wechseln Sie zu &quot;Beschaffung&quot; &gt; &quot;Angebotsanforderungen&quot; &gt; &quot;Alle Angebotsanforderungen&quot;.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="44">Klicken Sie auf &quot;Neu&quot;.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="45">Wählen Sie im Feld &quot;Ausschreibungstyp&quot; den Ausschreibungstyp aus, den Sie gerade erstellt haben.
*</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="47">Klicken Sie auf &quot;OK&quot;.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="48">Klicken Sie auf &quot;Bewertungskriterien&quot;.
<ul sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="49">
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="49">Die Bewertungskriterien, die angezeigt werden, sind diejenigen von der Bewertungsmethode, die Sie dem Ausschreibungstyp zugeordnet haben. Auf dieser Seite können Sie auswählen, Kriterien hinzuzufügen oder zu löschen. Es ist auch möglich, neue Kriterien hinzuzufügen, indem Sie diese aus anderen Bewertungsmethoden kopieren.</li>
</ul>
</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="50">Klicken Sie auf &quot;Kriterien kopieren&quot;.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="51">Geben Sie im Feld &quot;Bewertungsmethode&quot; einen Wert ein, oder wählen Sie einen Wert aus.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="52">Klicken Sie auf &quot;OK&quot;.</li>
<li sourcefile="articles_de/supply-chain/procurement/tasks/create-solicitation-types-scoring-criteria-rfqs.md" sourcestartlinenumber="53">Schließen Sie die Seite.</li>
</ol>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../../styles/main.js"></script>
  </body>
</html>
