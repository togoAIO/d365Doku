a   6  a   v     <  �  �  /  J  �  �     4  =  V  �        *  F    -     v   FileAndType�     �{"baseDir":"C:/D365-Operations/en-US/articles","file":"human-resources/hr-leave-and-absence-analytics.md","type":"article","sourceDir":"","destinationDir":""}   <  OriginalFileAndType�   �  �{"baseDir":"C:/D365-Operations/en-US/articles","file":"human-resources/hr-leave-and-absence-analytics.md","type":"article","sourceDir":"","destinationDir":""}   �  Key=   /  3~/human-resources/hr-leave-and-absence-analytics.md   J  LocalPathFromRoot;   �  1human-resources/hr-leave-and-absence-analytics.md   �  LinkToFiles      �  �  9   �  /~/human-resources/hr-leave-and-absence-plans.md<      2~/human-resources/hr-leave-and-absence-overview.md   4  
LinkToUids	   =     V  FileLinkSources�  �  �{"~/human-resources/hr-leave-and-absence-plans.md":[{"Target":"~/human-resources/hr-leave-and-absence-plans.md","SourceFile":"human-resources/hr-leave-and-absence-analytics.md","LineNumber":51}],"~/human-resources/hr-leave-and-absence-overview.md":[{"Target":"~/human-resources/hr-leave-and-absence-overview.md","SourceFile":"human-resources/hr-leave-and-absence-analytics.md","LineNumber":50}]}     UidLinkSources     {}     Uids   *  []   F  ManifestProperties�     �{"rawTitle":"<h1 id=\"view-analytics-for-leave-and-absence\" sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"32\">View analytics for leave and absence</h1>"}   -  DocumentType	   6     <$  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","conceptual":"\n<p sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"34\">Dynamics 365 Human Resources provides analytics to help give you insight into your organization's leave and absence trends.</p>\n<h2 id=\"view-leave-and-absence-analytics\" sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"36\">View Leave and absence analytics</h2>\n<ol sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"38\">\n<li sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"38\"><p sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"38\">In the <strong sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"38\">Leave and absence</strong> workspace, select the <strong sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"38\">Analytics</strong> tab.</p>\n</li>\n<li sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"40\"><p sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"40\">Choose one of the following views from the tabs along the bottom:</p>\n<ul sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"42\">\n<li sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"42\"><p sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"42\"><strong sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"42\">Leave and Absence Overview</strong> - View enrollment percentages and utilization rates for your leave plans, monthly accruals and balances, and time-off balances by manager.</p>\n</li>\n<li sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"44\"><p sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"44\"><strong sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"44\">Current Balance Analysis</strong> - View detailed information about leave balances and accruals.</p>\n</li>\n<li sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"46\"><p sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"46\"><strong sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"46\">Balance Trend Analysis</strong> - View trends in leave balances by month and by year, and view trends over the past 12 months.</p>\n</li>\n</ul>\n</li>\n</ol>\n<h2 id=\"see-also\" sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"48\">See also</h2>\n<ul sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"50\">\n<li sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"50\"><a href=\"~/human-resources/hr-leave-and-absence-overview.md\" sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"50\">Leave and absence overview</a></li>\n<li sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"51\"><a href=\"~/human-resources/hr-leave-and-absence-plans.md\" sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"51\">Create a leave and absence plan</a></li>\n</ul>\n","type":"Conceptual","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"articles/human-resources/hr-leave-and-absence-analytics.md","branch":"live","repo":"https://github.com/MicrosoftDocs/Dynamics-365-unified-Operations-public"},"startLine":0,"endLine":0,"isExternal":false},"path":"human-resources/hr-leave-and-absence-analytics.md","documentation":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"articles/human-resources/hr-leave-and-absence-analytics.md","branch":"live","repo":"https://github.com/MicrosoftDocs/Dynamics-365-unified-Operations-public"},"startLine":0,"endLine":0,"isExternal":false},"layout":"Conceptual","search.app":{"$type":"System.Object[], mscorlib","$values":["HumanResources"]},"feedback_github_repo":"MicrosoftDocs/dynamics-365-unified-operations-public","ms.search.scope":"Core, Operations, Human Resources, ShowInHelp","feedback_system":"GitHub","_norobots":true,"feedback_product_url":"https://ideas.dynamics.com","breadcrumb_path":"/dynamics365/ops-bc/toc.json","_docfxVersion":"2.56.6.0","titleSuffix":"Human Resources | Dynamics 365","_op_documentIdPathDepotMapping":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","dev-itpro/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsDevITPro"},"financials/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsFinancials"},"fin-and-ops/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsCore"},"retail/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsRetail"},"supply-chain/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsSCM"},"talent/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsHR"}},"extendBreadcrumb":"true","contributors_to_exclude":{"$type":"System.Object[], mscorlib","$values":["OpenLocalizationService","buck1ey","bishalgoswami"]},"searchScope":{"$type":"System.Object[], mscorlib","$values":["Dynamics 365","Unified Operations","Human Resources"]},"brand":"dyn-ops","uhfHeaderId":"MSDocsHeader-Dynamics365","_noindex":true,"_systemKeys":{"$type":"System.String[], mscorlib","$values":["conceptual","type","source","path","documentation","title","rawTitle","wordCount"]},"rawTitle":"<h1 id=\"view-analytics-for-leave-and-absence\" sourcefile=\"human-resources/hr-leave-and-absence-analytics.md\" sourcestartlinenumber=\"32\">View analytics for leave and absence</h1>","ms.custom":7521,"title":"View analytics for leave and absence","ms.dyn365.ops.version":"Human Resources","ms.search.region":"Global","ms.assetid":null,"author":"andreabichsel","description":"View leave analytics, accruals and balances, and balance trends in Dynamics 365 Human Resources.","ms.author":"anbichse","audience":"Application User","manager":"AnnBe","ms.search.validFrom":"2020-02-03","ms.topic":"article","ms.search.form":"LeavePlanFormPart, LeaveAbsenceWorkspace","ms.service":"dynamics-human-resources","ms.date":"02/03/2020","ms.technology":null,"ms.prod":null,"ms.reviewer":"anbichse"}�   �$  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","IsUserDefinedTitle":true,"XrefSpec":null}	   �$   