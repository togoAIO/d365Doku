a   �
  a   v   &  C  �     =  X  �  �  �  �      7	  O	  [	  i	  u	  �	  l
  �
     v   FileAndType�   &  �{"baseDir":"C:/D365-Operations/OwnDocu/d365Doku_D365","file":"articles/commerce/experimentation-connect-edit.md","type":"article","sourceDir":"","destinationDir":""}   C  OriginalFileAndType�   �  �{"baseDir":"C:/D365-Operations/OwnDocu/d365Doku_D365","file":"articles/commerce/experimentation-connect-edit.md","type":"article","sourceDir":"","destinationDir":""}      Key=   =  3~/articles/commerce/experimentation-connect-edit.md   X  LocalPathFromRoot;   �  1articles/commerce/experimentation-connect-edit.md   �  LinkToFiles   �  �  	  ?    �  D   	  :~/articles/commerce/media/experimentation_connect_edit.svg6   ?  ,~/articles/commerce/experimentation-setup.md@     6~/articles/commerce/experimentation-preview-publish.md/   �  %~/articles/commerce/publish-groups.md9   �  /~/articles/commerce/experimentation-overview.md   �  
LinkToUids	          FileLinkSources  7	  �
{"~/articles/commerce/media/experimentation_connect_edit.svg":[{"Target":"~/articles/commerce/media/experimentation_connect_edit.svg","Anchor":"#lightbox","SourceFile":"articles/commerce/experimentation-connect-edit.md","LineNumber":37},{"Target":"~/articles/commerce/media/experimentation_connect_edit.svg","SourceFile":"articles/commerce/experimentation-connect-edit.md","LineNumber":37}],"~/articles/commerce/experimentation-setup.md":[{"Target":"~/articles/commerce/experimentation-setup.md","SourceFile":"articles/commerce/experimentation-connect-edit.md","LineNumber":39},{"Target":"~/articles/commerce/experimentation-setup.md","SourceFile":"articles/commerce/experimentation-connect-edit.md","LineNumber":96}],"~/articles/commerce/experimentation-preview-publish.md":[{"Target":"~/articles/commerce/experimentation-preview-publish.md","SourceFile":"articles/commerce/experimentation-connect-edit.md","LineNumber":100}],"~/articles/commerce/publish-groups.md":[{"Target":"~/articles/commerce/publish-groups.md","SourceFile":"articles/commerce/experimentation-connect-edit.md","LineNumber":58}],"~/articles/commerce/experimentation-overview.md":[{"Target":"~/articles/commerce/experimentation-overview.md","SourceFile":"articles/commerce/experimentation-connect-edit.md","LineNumber":74}]}   O	  UidLinkSources   [	  {}   i	  Uids   u	  []   �	  ManifestProperties�   l
  �{"rawTitle":"<h1 id=\"connect-an-experiment-and-edit-variations\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"31\">Connect an experiment and edit variations</h1>"}   �
  DocumentType	   �
   �>  3I  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","conceptual":"\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"33\">This topic describes how to connect your experiment in Commerce and make changes to your variations so that they align with your hypothesis.</p>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"35\">The following diagram shows all of the steps involved in setting up and running an experiment on an e-Commerce website in Dynamics 365 Commerce. Additional steps are covered in separate topics.</p>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"37\"><a href=\"~/articles/commerce/media/experimentation_connect_edit.svg#lightbox\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"37\"> <img src=\"~/articles/commerce/media/experimentation_connect_edit.svg\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"37\" alt=\"Experimentation user journey - Connect &amp; Edit\"> </a></p>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"39\">After you've <a href=\"~/articles/commerce/experimentation-setup.md\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"39\">set up your experiment</a> in a third-party service, you'll connect the experiment in Dynamics 365 Commerce and edit the experiment variations.</p>\n<h2 id=\"planning-considerations\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"41\">Planning considerations</h2>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"43\">Before you connect your experiment in Commerce, you'll need to make some decisions that impact the way Commerce manages your content.</p>\n<h3 id=\"determine-the-scope-of-your-experiment\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"45\">Determine the scope of your experiment</h3>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"46\">When you connect an experiment, you are prompted to define the scope of the experiment. Experiments are defined as <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"46\">partial</strong> scope or <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"46\">entire</strong> scope.</p>\n<ul sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"47\">\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"47\">Choose <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"47\">partial</strong> if you want to conduct an experiment on a specific portion of a page. If you select this option, you must identify which modules are included in the experiment. Changes that are made to parts of the default page or fragment that aren't related to the experiment are automatically synchronized across variations.</li>\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"48\">Choose <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"48\">entire</strong> if you want to conduct an experiment on an entire page or fragment. Separate copies of the default page or fragment are created. You won't have to select which modules are included in the experiment because the whole editing surface is available to change. You can add, delete, or re-order modules as needed. However, if any changes are made to the default page or fragment that the experiment is associated with, those changes have to be manually synchronized across all variations.</li>\n</ul>\n<!-- not to editors, we're adding an image here to illustrate the difference. it will help.) -->\n<div class=\"NOTE\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"52\">\n<h5>Note</h5>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"53\">If you associate your experiment with a page that uses a layout, you can only scope the experiment as <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"53\">entire</strong>.</p>\n</div>\n<h3 id=\"decide-if-you-want-to-schedule-when-your-experiment-is-published\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"55\">Decide if you want to schedule when your experiment is published</h3>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"56\">If you want to schedule when your experiment is published to your live site, make sure the content you want to associate with the experiment is available in a publish group <em sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"56\">before</em> you connect the experiment.</p>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"58\">For more information about publish groups, refer to <a href=\"~/articles/commerce/publish-groups.md\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"58\">Work with publish groups</a>.</p>\n<h2 id=\"connect-your-experiment\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"61\">Connect your experiment</h2>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"62\">To connect your experiment, you'll launch the <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"62\">Connect experiment</strong> wizard. The wizard walks you through the steps required to connect your experiment. When you complete the wizard, your experiment is connected and variations are created and ready to be edited.</p>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"64\">To get started connecting your experiment in Commerce site builder, follow these steps.</p>\n<ol sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"66\">\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"66\"><p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"66\">To launch the <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"66\">Connect experiment</strong> wizard, select <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"66\">Experiments</strong> in the left navigation pane, and then select <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"66\">Connect</strong>. Alternatively, you can access the wizard from a page or fragment editor by editing it and selecting <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"66\">Connect experiment</strong> on the command bar.</p>\n<div class=\"NOTE\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"68\">\n<h5>Note</h5>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"69\">A page can only be connected to one experiment at a time. To connect a page to a different experiment, first delete the experiment that the page is currently connected to.</p>\n</div>\n</li>\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"71\"><p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"71\">Choose the page or fragment you want to run your experiment on.</p>\n</li>\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"72\"><p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"72\">Set the experimentation scope to <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"72\">partial</strong> or <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"72\">entire</strong>, based on the choice you made in the <a href=\"#determine-the-scope-of-your-experiment\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"72\">Determine the scope of your experiment</a> section above.</p>\n<div class=\"NOTE\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"73\">\n<h5>Note</h5>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"74\">The <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"74\">Experiment on pages or fragments</strong> feature flag must be enabled if you want to experiment on a full page or fragment. Refer to the <a href=\"~/articles/commerce/experimentation-overview.md\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"74\">Experimentation in Dynamics 365 Commerce</a> topic for more information.</p>\n</div>\n</li>\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"76\"><p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"76\">In the final step of the wizard, select <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"76\">Generate variations and exit wizard</strong>. Variations are created for the experiment.</p>\n</li>\n</ol>\n<h2 id=\"edit-your-variations\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"78\">Edit your variations</h2>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"79\">When you exit the wizard, variations are created for you.</p>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"81\">Next, you'll edit the variations so they reflect the choices that you need to verify in the experiment hypothesis. Choose one of following procedures that corresponds to the scope you chose for your experiment in the <a href=\"#determine-the-scope-of-your-experiment\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"81\">Determine the scope of your experiment</a> section above.</p>\n<h3 id=\"edit-variations-for-experiments-with-partial-scope\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"83\">Edit variations for experiments with partial scope</h3>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"84\">Follow these steps if you defined the scope of your experiment as <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"84\">partial</strong> in the <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"84\">Connect experiment</strong> wizard.</p>\n<ol sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"86\">\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"86\">In editor view, use the variations drop-down menu below the command bar to edit each variation based on your original hypothesis. You may also want to establish a control or base variation by leaving one of the variations unchanged.</li>\n<li sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"87\">Select the module to be experimented on, select the ellipsis (...), and then select <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"87\">Add to experiment</strong>.</li>\n</ol>\n<h3 id=\"edit-variations-for-experiments-with-entire-scope\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"89\">Edit variations for experiments with entire scope</h3>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"90\">If you defined the scope of your experiment as <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"90\">entire</strong> in the <strong sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"90\">Connect experiment</strong> wizard, while in editor view, use the variations drop-down menu below the command bar to edit each variation based on your original hypothesis.</p>\n<div class=\"NOTE\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"92\">\n<h5>Note</h5>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"93\">In either case, you may also want to establish a control or base variation by leaving one of the variations unchanged.</p>\n</div>\n<h2 id=\"previous-step\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"95\">Previous step</h2>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"96\"><a href=\"~/articles/commerce/experimentation-setup.md\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"96\">Set up an experiment</a></p>\n<h2 id=\"next-step\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"99\">Next step</h2>\n<p sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"100\"><a href=\"~/articles/commerce/experimentation-preview-publish.md\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"100\">Preview and publish an experiment</a></p>\n","type":"Conceptual","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"articles/commerce/experimentation-connect-edit.md","branch":"main","repo":"https://github.com/togoAIO/d365Doku.git"},"startLine":0,"endLine":0,"isExternal":false},"path":"articles/commerce/experimentation-connect-edit.md","documentation":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"articles/commerce/experimentation-connect-edit.md","branch":"main","repo":"https://github.com/togoAIO/d365Doku.git"},"startLine":0,"endLine":0,"isExternal":false},"_enableSearch":"true","_docfxVersion":"2.56.6.0","_appTitle":"WIKA Documentation","_systemKeys":{"$type":"System.String[], mscorlib","$values":["conceptual","type","source","path","documentation","title","rawTitle","wordCount"]},"rawTitle":"<h1 id=\"connect-an-experiment-and-edit-variations\" sourcefile=\"articles/commerce/experimentation-connect-edit.md\" sourcestartlinenumber=\"31\">Connect an experiment and edit variations</h1>","ms.custom":null,"title":"Connect an experiment and edit variations","ms.dyn365.ops.version":"AX 10.0.13","ms.search.region":"global","ms.assetid":null,"author":"sushma-rao","description":"This topic describes how to connect an experiment in a third-party service to Dynamics 365 Commerce, and how to edit variations for the experiment.","ms.author":"sushmar","audience":"Application User","manager":"AnnBe","ms.search.validFrom":"2020-09-30","ms.topic":"article","ms.service":"dynamics-365-retail","ms.search.industry":"Retail","ms.date":"10/21/2020","ms.technology":null,"ms.prod":null,"ms.reviewer":"josaw"}�   �I  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","IsUserDefinedTitle":true,"XrefSpec":null}	   �I   