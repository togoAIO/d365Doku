a   �	  a   v   2  O      h  �  �  �    3  <  U  -  E  Q  _  k  �  c	  y	     v   FileAndType�   2  �{"baseDir":"C:/D365-Operations/en-US/articles","file":"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","type":"article","sourceDir":"","destinationDir":""}   O  OriginalFileAndType�     �{"baseDir":"C:/D365-Operations/en-US/articles","file":"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","type":"article","sourceDir":"","destinationDir":""}     KeyP   h  F~/finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md   �  LocalPathFromRootN   �  Dfinance/localizations/apac-ind-GST-purchase-from-composite-dealer.md   �  LinkToFiles     �  G  �  �  H   G  >~/finance/localizations/media/Annotation-2019-05-16-100656.pngH   �  >~/finance/localizations/media/Annotation-2019-05-16-101138.pngH   �  >~/finance/localizations/media/Annotation-2019-05-16-101054.pngH     >~/finance/localizations/media/Annotation-2019-05-16-101246.png   3  
LinkToUids	   <     U  FileLinkSources�  -  �{"~/finance/localizations/media/Annotation-2019-05-16-100656.png":[{"Target":"~/finance/localizations/media/Annotation-2019-05-16-100656.png","SourceFile":"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","LineNumber":62}],"~/finance/localizations/media/Annotation-2019-05-16-101138.png":[{"Target":"~/finance/localizations/media/Annotation-2019-05-16-101138.png","SourceFile":"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","LineNumber":43}],"~/finance/localizations/media/Annotation-2019-05-16-101054.png":[{"Target":"~/finance/localizations/media/Annotation-2019-05-16-101054.png","SourceFile":"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","LineNumber":39}],"~/finance/localizations/media/Annotation-2019-05-16-101246.png":[{"Target":"~/finance/localizations/media/Annotation-2019-05-16-101246.png","SourceFile":"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","LineNumber":47}]}   E  UidLinkSources   Q  {}   _  Uids   k  []   �  ManifestProperties�   c	  �{"rawTitle":"<h1 id=\"purchases-from-composite-dealers\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"30\">Purchases from composite dealers</h1>"}   y	  DocumentType	   �	    *  �3  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","conceptual":"\n\n<ol sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"34\">\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"34\"><p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"34\">Go to <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"34\">Accounts payable</strong> &gt; <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"34\">Invoice</strong> &gt; <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"34\">Invoice journals</strong>.</p>\n</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"35\"><p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"35\">Create a journal, and then select <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"35\">Lines</strong>.</p>\n</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"36\"><p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"36\">Create a purchase transaction for a composite vendor, and save the record.</p>\n</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"37\"><p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"37\">Select <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"37\">Tax information</strong>.</p>\n<p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"39\"><img src=\"~/finance/localizations/media/Annotation-2019-05-16-101054.png\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"39\" alt=\"Tax information dialog box\"></p>\n</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"41\"><p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"41\">On the <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"41\">GST</strong> FastTab, in the <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"41\">HSN codes</strong> field, select a value.</p>\n<p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"43\"><img src=\"~/finance/localizations/media/Annotation-2019-05-16-101138.png\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"43\" alt=\"GST FastTab\"></p>\n</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"45\"><p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"45\">On the <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"45\">Vendor tax information</strong> FastTab, verify the information.</p>\n<p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"47\"><img src=\"~/finance/localizations/media/Annotation-2019-05-16-101246.png\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"47\" alt=\"Vendor tax information FastTab\"></p>\n</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"49\"><p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"49\">Select <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"49\">OK</strong>.</p>\n</li>\n</ol>\n<h2 id=\"validate-the-tax-details\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"51\">Validate the tax details</h2>\n<ol sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"53\">\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"53\">Select <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"53\">Tax document</strong>.</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"54\">Select <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"54\">Close</strong>.</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"55\">Select <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"55\">Post</strong> &gt; <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"55\">Post</strong> to post the journal.</li>\n<li sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"56\">Close the message that you receive.</li>\n</ol>\n<h2 id=\"validate-a-voucher\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"58\">Validate a voucher</h2>\n<p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"60\">To validate a voucher, select <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"60\">Inquiries</strong> &gt; <strong sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"60\">Voucher</strong>.</p>\n<p sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"62\"><img src=\"~/finance/localizations/media/Annotation-2019-05-16-100656.png\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"62\" alt=\"Example\"></p>\n","type":"Conceptual","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"articles/finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","branch":"live","repo":"https://github.com/MicrosoftDocs/Dynamics-365-unified-Operations-public"},"startLine":0,"endLine":0,"isExternal":false},"path":"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","documentation":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"articles/finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md","branch":"live","repo":"https://github.com/MicrosoftDocs/Dynamics-365-unified-Operations-public"},"startLine":0,"endLine":0,"isExternal":false},"layout":"Conceptual","search.app":{"$type":"System.Object[], mscorlib","$values":["Finance"]},"feedback_github_repo":"MicrosoftDocs/dynamics-365-unified-operations-public","ms.search.scope":"Core, Operations, Finance","feedback_system":"GitHub","_norobots":true,"feedback_product_url":"https://ideas.dynamics.com","breadcrumb_path":"/dynamics365/ops-bc/toc.json","_docfxVersion":"2.56.6.0","titleSuffix":"Finance | Dynamics 365","_op_documentIdPathDepotMapping":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","dev-itpro/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsDevITPro"},"financials/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsFinancials"},"fin-and-ops/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsCore"},"retail/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsRetail"},"supply-chain/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsSCM"},"talent/":{"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","folder_relative_path_in_docset":".","depot_name":"MSDN.d365OpsHR"}},"extendBreadcrumb":"true","contributors_to_exclude":{"$type":"System.Object[], mscorlib","$values":["OpenLocalizationService","buck1ey","bishalgoswami"]},"searchScope":{"$type":"System.Object[], mscorlib","$values":["Dynamics 365","Unified Operations"]},"brand":"dyn-ops","uhfHeaderId":"MSDocsHeader-Dynamics365","_noindex":true,"_systemKeys":{"$type":"System.String[], mscorlib","$values":["conceptual","type","source","path","documentation","title","rawTitle","wordCount"]},"rawTitle":"<h1 id=\"purchases-from-composite-dealers\" sourcefile=\"finance/localizations/apac-ind-GST-purchase-from-composite-dealer.md\" sourcestartlinenumber=\"30\">Purchases from composite dealers</h1>","title":"Purchases from composite dealers","ms.dyn365.ops.version":"10.0.4","ms.search.region":"India","author":"EricWang","description":"This topic provides information about purchases that are made from a composite dealer.","ms.author":"kfend","audience":"Application User","manager":"RichardLuan","ms.search.validFrom":"2019-06-01","ms.topic":"article","ms.service":"dynamics-365-applications","ms.date":"06/04/2019","ms.technology":null,"ms.prod":null,"ms.reviewer":"kfend"}�   G4  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","IsUserDefinedTitle":true,"XrefSpec":null}	   P4   