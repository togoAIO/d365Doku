<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Liste der EB-Funktionen in der Typenumrechnungskategorie | WIKA Documentation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Liste der EB-Funktionen in der Typenumrechnungskategorie | WIKA Documentation ">
    <meta name="generator" content="docfx 2.56.6.0">
    
    <link rel="shortcut icon" href="../../../../microsoft-dynamics-crm-365-icon.ico">
    <link rel="stylesheet" href="../../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../../styles/main.css">
    <link href="https://fonts.googleapis.com/css?family=Roboto" rel="stylesheet"> 
    <meta property="docfx:navrel" content="../../../../toc.html">
    <meta property="docfx:tocrel" content="../../../commerce/TOC.html">
    
    <meta property="docfx:rel" content="../../../../">
    
  </head>  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../../index.html">
                <img id="logo" class="svg" src="../../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div class="container body-content">
        
        <div id="search-results">
          <div class="search-list">Search Results for <span></span></div>
          <div class="sr-items">
            <p><i class="glyphicon glyphicon-refresh index-loading"></i></p>
          </div>
          <ul id="pagination" data-first="First" data-prev="Previous" data-next="Next" data-last="Last"></ul>
        </div>
      </div>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="">
<h1 id="list-of-er-functions-in-the-type-conversion-category" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="27">Liste der EB-Funktionen in der Typenumrechnungskategorie</h1>

[!include[banner](../includes/banner.md)]
<p sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="31">Konvertierungsfunktionen für EB-Typen (elektronische Berichterstellung) können zum Konvertieren von Werten zwischen Typen verwendet werden. Dieses Thema enthält eine Zusammenfassung dieser Funktionen.</p>
<h2 id="type-conversion-functions" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="33">Funktionen zur Typenumrechnung</h2>
<table sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="35">
<thead>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="35">
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="35">Funktion</th>
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="35">Beschreibung</th>
</tr>
</thead>
<tbody>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="37">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="37"><a href="er-functions-conversion-int64value.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="37">Int64Value</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="37">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="37">Int64</em> zurück, der die angegebene Zeichenfolge darstellt.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="38">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="38"><a href="er-functions-conversion-intvalue.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="38">IntValue</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="38">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="38">Int</em> zurück, der die angegebene Zeichenfolge darstellt.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="39">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="39"><a href="er-functions-conversion-numbervalue.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="39">NumberValue</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="39">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="39">Real</em> zurück, der über den angegebenen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="39">String</em> konvertiert wird. Bei der Konvertierung werden die angegebenen Trennzeichen für Dezimal- und Zifferngruppierungen berücksichtigt.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="40">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="40"><a href="er-functions-conversion-value.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="40">Wert</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="40">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="40">Real</em> zurück, der über den angegebenen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="40">String</em> konvertiert wird.</td>
</tr>
</tbody>
</table>
<h2 id="type-conversion-functions-in-the-date-and-time-category" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="42">Typenumrechnungsfunktionen in der Kategorie „Datum und Uhrzeit“</h2>
<p sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="44">Die folgende Tabelle beschreibt die Typenumrechnungsfunktionen in der <a href="er-functions-category-datetime.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="44">Kategorie „Datum und Uhrzeit“</a>.</p>
<table sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="46">
<thead>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="46">
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="46">Funktion</th>
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="46">Beschreibung</th>
</tr>
</thead>
<tbody>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="48">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="48"><a href="er-functions-datetime-datetimevalue.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="48">DateTimeValue</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="48">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="48">DateTime</em> zurück, der über den vorgegebenen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="48">String</em> im speziellen Format und in der optional angegebenen Kultur in den Wert für Datum/Uhrzeit konvertiert wird.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="49">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="49"><a href="er-functions-datetime-datetodatetime.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="49">DateToDateTime</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="49">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="49">DateTime</em> zurück, der über den vorgegebenen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="49">Date</em> in einen Wert für Datum/Uhrzeit in der Koordinierten Weltzeit (Greenwich Mean Time [GMT]) konvertiert wird.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="50">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="50"><a href="er-functions-datetime-datevalue.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="50">DateValue</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="50">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="50">Date</em> zurück, der über den vorgegebenen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="50">String</em> im speziellen Format und in der optional angegebenen Kultur in den Wert für Datum konvertiert wird.</td>
</tr>
</tbody>
</table>
<h2 id="type-conversion-functions-in-the-list-category" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="52">Typenumrechnungsfunktionen in der Listenkategorie</h2>
<p sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="54">Die folgende Tabelle beschreibt die Typenumrechnungsfunktionen in der <a href="er-functions-category-list.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="54">Listenkategorie</a>.</p>
<table sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="56">
<thead>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="56">
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="56">Funktion</th>
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="56">Beschreibung</th>
</tr>
</thead>
<tbody>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="58">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="58"><a href="er-functions-list-list.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="58">Liste</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="58">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="58">Datensatzliste</em> als neue Liste zurück, die anhand der angegebenen Argumente des Typs <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="58">Container (Datensatz)</em> erstellt wird.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="59">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="59"><a href="er-functions-list-listoffields.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="59">ListOfFields</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="59">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="59">Datensatzliste</em> zurück, der basierend auf der Struktur des angegebenen Arguments des Typs <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="59">Aufzählung</em> oder <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="59">Container (Datensatz)</em> erstellt wird.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="60">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="60"><a href="er-functions-list-split.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="60">Teilen</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="60">Diese Funktion teilt den angegebenen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="60">String</em> in Teilzeichenfolgen auf und gibt das Ergebnis als neuen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="60">Datensatzliste</em> zurück.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="61">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="61"><a href="er-functions-list-stringjoin.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="61">StringJoin</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="61">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="61">String</em> zurück, der aus verketteten Werten des angegebenen Feldes aus dem angegebenen Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="61">Datensatzliste</em> besteht. Die Werte können durch das angegebene Trennzeichen getrennt werden.</td>
</tr>
</tbody>
</table>
<h2 id="type-conversion-functions-in-the-text-category" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="63">Typenumrechnungsfunktionen in der Textkategorie</h2>
<p sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="65">Die folgende Tabelle beschreibt die Typenumrechnungsfunktionen in der <a href="er-functions-category-text.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="65">Textkategorie</a>.</p>
<table sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="67">
<thead>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="67">
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="67">Funktion</th>
<th sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="67">Beschreibung</th>
</tr>
</thead>
<tbody>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="69">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="69"><a href="er-functions-text-char.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="69">Char</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="69">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="69">String</em> zurück, der ein einzelnes Zeichen darstellt, auf das durch die angegebene Unicode-Nummer verwiesen wird.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="70">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="70"><a href="er-functions-text-guidvalue.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="70">GuidValue</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="70">Diese Funktion konvertiert die angegebene Eingabe des Datentyps <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="70">String</em> in ein Datenelement des Typs <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="70">GUID</em>.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="71">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="71"><a href="er-functions-text-numberformat.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="71">NumberFormat</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="71">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="71">String</em> zurück, der eine angegebene Zahl im angegebenen Format und in einer optional angegebenen Kultur darstellt.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="72">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="72"><a href="er-functions-text-qrcode.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="72">QrCode</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="72">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="72">Container</em> zurück, der das QR-Code-Bild (Quick Response Code) für die angegebene Zeichenfolge im Binärformat darstellt.</td>
</tr>
<tr sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="73">
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="73"><a href="er-functions-text-text.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="73">Text</a></td>
<td sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="73">Diese Funktion gibt den Wert <em sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="73">String</em> zurück, der die angegebene Zahl darstellt, nachdem sie in eine Textzeichenfolge konvertiert wurde, die gemäß den Servergebietsschemaeinstellungen der aktuellen Anwendungsinstanz formatiert ist.</td>
</tr>
</tbody>
</table>
<h2 id="additional-resources" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="75">Zusätzliche Ressourcen</h2>
<p sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="77"><a href="general-electronic-reporting.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="77">Überblick über die elektronische Berichterstellung</a></p>
<p sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="79"><a href="general-electronic-reporting-formula-designer.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="79">Formeldesigner in der elektronischen Berichterstellung</a></p>
<p sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="81"><a href="er-formula-language.html" sourcefile="articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md" sourcestartlinenumber="81">Formelsprache in der elektronischen Berichterstellung</a></p>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                  <li>
                    <a href="https://github.com/togoAIO/d365Doku/blob/main/articles_de/fin-ops-core/dev-itpro/analytics/er-functions-category-type-conversion.md/#L1" class="contribution-link">Improve this Doc</a>
                  </li>
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../../styles/main.js"></script>
  </body>
</html>
