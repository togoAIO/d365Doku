<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>What's new or changed in Dynamics 365 Supply Chain Management 10.0.7 (January 2020) | WIKA Documentation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="What's new or changed in Dynamics 365 Supply Chain Management 10.0.7 (January 2020) | WIKA Documentation ">
    <meta name="generator" content="docfx 2.56.6.0">
    
    <link rel="shortcut icon" href="../../../microsoft-dynamics-crm-365-icon.ico">
    <link rel="stylesheet" href="../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../styles/main.css">
    <link href="https://fonts.googleapis.com/css?family=Roboto" rel="stylesheet"> 
    <meta property="docfx:navrel" content="../../../toc.html">
    <meta property="docfx:tocrel" content="../toc.html">
    
    
    
  </head>  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../index.html">
                <img id="logo" class="svg" src="../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="">
<h1 id="whats-new-or-changed-in-dynamics-365-supply-chain-management-1007-january-2020" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="32">What's new or changed in Dynamics 365 Supply Chain Management 10.0.7 (January 2020)</h1>


<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="37">This topic describes features that are either new or changed in Microsoft Dynamics 365 Supply Chain Management 10.0.7. This version has a build number of 10.0.283, and is available as follows:</p>
<ul sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="39">
<li sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="39">Preview release is in October 2019.</li>
<li sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="40">General availability (self-update) is in November 2019.</li>
<li sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="41">Auto-update is in January 2020.</li>
</ul>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="43">For more information about version 10.0.7, see <a href="whats-new-scm-10-0-7.html#additional-resources" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="43">Additional resources</a>.</p>
<h2 id="feature-management-enhancements" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="45">Feature management enhancements</h2>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="46">Feature management now allows you to enable all new features by default, require confirmation to enable a feature, and enable all features that have not already been enabled.</p>
<h2 id="additional-resources" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="50">Additional resources</h2>
<h3 id="bug-fixes" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="52">Bug fixes</h3>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="53">For information about the bug fixes included in each of the updates that are part of 10.0.7, sign in to Lifecycle Services (LCS) and view the <a href="https://fix.lcs.dynamics.com/Issue/Details?kb=4528173&amp;bugId=386529&amp;dbType=3&amp;qc=d6f5cd3ead06907477eae511043a52c1d4290a12bf52374dd55faf0d28ae732e" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="53">KB article</a>.</p>
<h3 id="platform-update-31" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="55">Platform update 31</h3>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="56">Microsoft Dynamics 365 Supply Chain Management 10.0.7 includes Platform update 31. To learn more about Platform update 31, see <a href="https://docs.wika.com/en-us/dynamics365/supply-chain/fin-ops-core/dev-itpro/get-started/whats-new-platform-update-31" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="56">What's new or changed in Platform update 31 (This is an external linThis link was changed due to HTMLfromRepoGenerator)</a>.</p>
<h3 id="dynamics-365-2019-release-wave-2-plan" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="58">Dynamics 365: 2019 release wave 2 plan</h3>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="59">Wondering about upcoming and recently released capabilities in any of our business apps or platform?</p>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="61">Check out the <a href="https://docs.microsoft.com/dynamics365-release-plan/2019wave2/" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="61">Dynamics 365: 2019 release wave 2 plan</a>. We've captured all the details, end to end, top to bottom, in a single document that you can use for planning.</p>
<h3 id="removed-and-deprecated-supply-chain-management-features" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="63">Removed and deprecated Supply Chain Management features</h3>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="65">The <a href="removed-deprecated-features-scm-updates.html" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="65">Removed or deprecated features in Dynamics 365 Supply Chain Management</a> topic describes features that have been or are scheduled to be removed or deprecated for Supply Chain Management.</p>
<ul sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="67">
<li sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="67">A <em sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="67">removed</em> feature is no longer available in the product.</li>
<li sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="68">A <em sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="68">deprecated</em> feature is not in active development and may be removed in a future update.</li>
</ul>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="70">Before any feature is removed from the product, the deprecation notice will be announced in the <a href="removed-deprecated-features-scm-updates.html" sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="70">Removed or deprecated features in Dynamics 365 Supply Chain Management</a> topic 12 months prior to the removal.</p>
<p sourcefile="articles/supply-chain/get-started/whats-new-scm-10-0-7.md" sourcestartlinenumber="72">For breaking changes that only affect compilation time, but are binary compatible with sandbox and production environments, the deprecation time will be less than 12 months. Typically, these are functional updates that need to be made to the compiler.</p>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../styles/main.js"></script>
  </body>
</html>
