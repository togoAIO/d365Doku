<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>E-Mail-Vorlagen verwalten | WIKA Documentation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="E-Mail-Vorlagen verwalten | WIKA Documentation ">
    <meta name="generator" content="docfx 2.56.6.0">
    
    <link rel="shortcut icon" href="../../../../../microsoft-dynamics-crm-365-icon.ico">
    <link rel="stylesheet" href="../../../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../../../styles/main.css">
    <link href="https://fonts.googleapis.com/css?family=Roboto" rel="stylesheet"> 
    <meta property="docfx:navrel" content="../../../../../toc.html">
    <meta property="docfx:tocrel" content="../../../../toc.html">
    
    
    
  </head>  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../../../index.html">
                <img id="logo" class="svg" src="../../../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="">
<h1 id="manage-email-templates" sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="25">E-Mail-Vorlagen verwalten</h1>

<div class="IMPORTANT" sourcefile="ProcessDoku/00_Basics/MS_Content/includes/banner.md" sourcestartlinenumber="1">
<h5>Important</h5>
</div>
<p sourcefile="ProcessDoku/00_Basics/MS_Content/includes/banner.md" sourcestartlinenumber="2">Diese Dokumentation ist teilweise von Microsoft verfasst und wurde nicht auf Vollständigkeit geprüft. Wenn informationen fehlen oder ein weiteres Kapitel hinzugefügt werden soll bitte eine Mail an das <a href="mailto:tobias.goldhammer@wika.com"></a> Dokumentations Team schreiben.</p>

<p sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="29">Sie können Informationen aus der Datenbank Ihrer Organisation in die Lesezeichen in einem neuen Dokument übertragen und in Vorlagen verwenden, die Sie bei der Kommunikation mit Bewerbern und Kandidaten unterstützen. Hierfür muss eine Vorlage mit Standardtext und einigen Lesezeichen an den Positionen erstellt werden, an denen die Systemdaten eingefügt werden sollen. So können Sie z. B. Adresse und Kontaktinformationen für einen Bewerber in ein Microsoft Word-Dokument einfügen, das Sie bei der Kommunikation mit diesem Bewerber verwenden können. Das Demodatenunternehmen, das verwendet wird, um diese Prozedur zu erstellen, ist USMF.</p>
<h2 id="select-which-bookmarks-to-use-in-your-email-templates" sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="32">Auswählen der Lesezeichen für die E-Mail-Vorlagen</h2>
<ol sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="33">
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="33">Gehen Sie im Navigationsbereich zu <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="33">Module &gt; Human Resources &gt; Recruitment &gt; Communication &gt; Application bookmarks</strong>.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="34">Suchen Sie in der Liste die gewünschten Korrespondenzaktivität, und wählen Sie sie aus.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="35">Wählen Sie <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="35">Bearbeiten</strong> aus.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="36">Wählen Sie die Felder aus, die Sie in einer E-Mail-Vorlage für die ausgewählte Korrespondenzaktivität verwenden möchten, und verschieben Sie sie in die Lesezeichenfelder.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="37">Schließen Sie die Seite.</li>
</ol>
<h2 id="create-an-email-template" sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="39">E-Mail-Vorlage erstellen</h2>
<ol sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="40">
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="40">Gehen Sie im Navigationsbereich zu <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="40">Module &gt; Personal &gt; Personalwesen &gt; Personalbeschaffung &gt; Kommunikation &gt; Vorlagen für Bewerbungs-E-Mails</strong>.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="41">Wählen Sie <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="41">Neu</strong> aus.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="42">Wählen Sie im Feld <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="42">Korrespondenzaktion</strong> <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="42">Interview</strong>. Wählen Sie die Korrespondenzaktivität aus, die Lesezeichen enthält, die für diese Art der E-Mail-Kommunikation verwendet wird.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="43">Geben Sie in das Feld <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="43">E-Mail-Vorlage</strong> einen Wert ein.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="44">Geben Sie in das Feld <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="44">Subjekt</strong> einen Wert ein.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="45">Geben Sie im Feld <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="45">Text</strong> einen Wert ein.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="46">Suchen Sie in der Liste das gewünschte Lesezeichenfeld, und wählen Sie es aus.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="47">Setzen Sie die Eingabe der E-Mail-Nachricht fort, und fügen Sie die Lesezeichenfelder an den gewünschten Positionen ein.</li>
<li sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="48">Wählen Sie <strong sourcefile="ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md" sourcestartlinenumber="48">Speichern</strong>.</li>
</ol>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../../../styles/main.js"></script>
  </body>
</html>
