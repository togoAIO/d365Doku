{
  "caution": "<p>Varning</p>",
  "classesInSubtitle": "Klasser",
  "constructorsInSubtitle": "Konstruktorer",
  "delegatesInSubtitle": "Delegeringar",
  "description": "Beskrivning",
  "eiisInSubtitle": "Explicita gränssnittsimplementeringar",
  "enumsInSubtitle": "Uppräkningar",
  "eventsInSubtitle": "Händelser",
  "examples": "Exempel",
  "exceptions": "Undantag",
  "extensionMethodsInSubtitle": "Tilläggsmetoder",
  "fieldsInSubtitle": "Fält",
  "fieldValue": "Fältvärde",
  "implements": "Implementeringar",
  "important": "<p>Viktigt</p>",
  "inheritance": "Arv",
  "inheritedMembers": "Ärvda medlemmar",
  "interfacesInSubtitle": "Gränssnitt",
  "inThisArticle": "I den här artikeln",
  "methodsInSubtitle": "Metoder",
  "name": "Namn",
  "namespace": "Namnområde",
  "note": "<p>Anteckning</p>",
  "operatorsInSubtitle": "Operatorer",
  "overrides": "Åsidosättningar",
  "parameters": "Parametrar",
  "propertiesInSubtitle": "Egenskaper",
  "propertyValue": "Egenskapsvärde",
  "remarks": "Kommentarer",
  "returns": "Returer",
  "seeAlso": "Se även",
  "structsInSubtitle": "Strukturer",
  "tip": "<p>Tips</p>",
  "type": "typ",
  "typeParameters": "Typparametrar",
  "warning": "<p>Varning</p>",

}